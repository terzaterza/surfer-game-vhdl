-- megafunction wizard: %ALTMEMMULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altmemmult 

-- ============================================================
-- File Name: hw_mult.vhd
-- Megafunction Name(s):
-- 			altmemmult
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altmemmult CBX_AUTO_BLACKBOX="ALL" COEFF_REPRESENTATION="UNSIGNED" COEFFICIENT0="79" DATA_REPRESENTATION="UNSIGNED" DEVICE_FAMILY="Cyclone III" MAX_CLOCK_CYCLES_PER_RESULT=1 RAM_BLOCK_TYPE="AUTO" TOTAL_LATENCY=2 WIDTH_C=8 WIDTH_D=8 WIDTH_R=16 clock data_in result
--VERSION_BEGIN 13.1 cbx_altaccumulate 2013:10:23:18:05:48:SJ cbx_altmemmult 2013:10:23:18:05:48:SJ cbx_altsyncram 2013:10:23:18:05:48:SJ cbx_cycloneii 2013:10:23:18:05:48:SJ cbx_lpm_add_sub 2013:10:23:18:05:48:SJ cbx_lpm_compare 2013:10:23:18:05:48:SJ cbx_lpm_counter 2013:10:23:18:05:48:SJ cbx_lpm_decode 2013:10:23:18:05:48:SJ cbx_lpm_mux 2013:10:23:18:05:48:SJ cbx_mgl 2013:10:23:18:06:54:SJ cbx_stratix 2013:10:23:18:05:48:SJ cbx_stratixii 2013:10:23:18:05:48:SJ cbx_stratixiii 2013:10:23:18:05:48:SJ cbx_stratixv 2013:10:23:18:05:48:SJ cbx_util_mgl 2013:10:23:18:05:48:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

--synthesis_resources = altsyncram 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  hw_mult_altmemmult_odo IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data_in	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 result_valid	:	OUT  STD_LOGIC
	 ); 
 END hw_mult_altmemmult_odo;

 ARCHITECTURE RTL OF hw_mult_altmemmult_odo IS

	 SIGNAL  wire_altsyncram1_q_a	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ECC_PIPELINE_STAGE_ENABLED	:	STRING := "FALSE";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTH_ECCSTATUS	:	NATURAL := 3;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone III";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(WIDTH_ECCSTATUS-1 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	result <= ( wire_altsyncram1_q_a(15 DOWNTO 0));
	result_valid <= '0';
	altsyncram1 :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "hw_mult.hex",
		OPERATION_MODE => "ROM",
		OUTDATA_REG_A => "CLOCK0",
		RAM_BLOCK_TYPE => "AUTO",
		WIDTH_A => 16,
		WIDTHAD_A => 8,
		INTENDED_DEVICE_FAMILY => "Cyclone III"
	  )
	  PORT MAP ( 
		address_a => data_in(7 DOWNTO 0),
		clock0 => clock,
		q_a => wire_altsyncram1_q_a
	  );

 END RTL; --hw_mult_altmemmult_odo
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY hw_mult IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data_in		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END hw_mult;


ARCHITECTURE RTL OF hw_mult IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT hw_mult_altmemmult_odo
	PORT (
			clock	: IN STD_LOGIC ;
			data_in	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(15 DOWNTO 0);

	hw_mult_altmemmult_odo_component : hw_mult_altmemmult_odo
	PORT MAP (
		clock => clock,
		data_in => data_in,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: COEFFICIENT0 STRING "79"
-- Retrieval info: PRIVATE: COEFF_REPRESENTATION_COMBO STRING "UNSIGNED"
-- Retrieval info: PRIVATE: COUNT_C_COMBO STRING "8"
-- Retrieval info: PRIVATE: COUNT_D_COMBO STRING "8"
-- Retrieval info: PRIVATE: DATA_REPRESENTATION_COMBO STRING "UNSIGNED"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: LOADABLE_COEFF STRING "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: SCLR_CHECK STRING "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: COEFFICIENT0 STRING "79"
-- Retrieval info: CONSTANT: COEFF_REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: DATA_REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: CONSTANT: MAX_CLOCK_CYCLES_PER_RESULT NUMERIC "1"
-- Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "AUTO"
-- Retrieval info: CONSTANT: TOTAL_LATENCY NUMERIC "2"
-- Retrieval info: CONSTANT: WIDTH_C NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_D NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_R NUMERIC "16"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_in 0 0 8 0 INPUT NODEFVAL "data_in[7..0]"
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL "result[15..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_in 0 0 8 0 data_in 0 0 8 0
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL hw_mult.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL hw_mult.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL hw_mult.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL hw_mult.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL hw_mult_inst.vhd FALSE
